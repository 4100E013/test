module test(in,out);

input in;
output reg ouy;

endmodule
